	module lights_off(sw, lights, clk, btn_fix, btn_rand, segment_led_1, segment_led_2);

	// control by switches
	input [9:0] sw;
	
	// stores the last status of the switches (helping the monitor of changes)
	reg [9:0] last = 10'b0000000000;
	
	// 50Mhz clock, pre-defined quiz, random quiz
	input clk, btn_fix, btn_rand;
	
	// indicate the current pre-defined quiz num
	reg fix_last = 0;
	
	// start count down if == 1
	reg start = 0;
	
	// cnt is the seconds ([7:4]=tens-dig, [3:0]=units_dig)
	reg [7:0] cnt;
	initial
	begin
		cnt[7:4] = 4'd0;
		cnt[3:0] = 4'd0;
	end
	
	// monitors if switches change on every posedge (true/false)
	reg [9:0] change = 10'b0000000000;
	
	// simulates a random value, increments on every posedge(50Mhz)
	reg [9:0] rd = 10'b0000000000;
	
	//increments on every posedge (50Mhz)(stablize the result)
	reg [23:0] fr; 
	
	// increments on every posedge (only coundown on 25-bit-one)
	reg [25:0] cd_fr;
	
	// connected to the led lights
	output reg [9:0] lights = 10'b0000000000;
	
	// parameter for xor operation (change state of specific lights)
	parameter [9:0] 
		c9 = 10'b1100000000,
		c8 = 10'b1110000000,
		c7 = 10'b0111000000,
		c6 = 10'b0011100000,
		c5 = 10'b0001110000,
		c4 = 10'b0000111000,
		c3 = 10'b0000011100,
		c2 = 10'b0000001110,
		c1 = 10'b0000000111,
		c0 = 10'b0000000011;
	
	// question number (0~4)
	reg [1:0] q_num = 0;
	
	// determine whether button is pressed (true/false)
	// change to next fixed question if true
	reg q_change = 0;
	
	// the pre-defined quizzes
	reg [9:0] q [3:0];
	initial
	begin
		q[0] = c0 ^ c1 ^ c2 ^ c3 ^ c4 ^ c5 ^ c6 ^ c7 ^ c8 ^ c9;	// answer: all
		q[1] = c0 ^ c2 ^ c3 ^ c5 ^ c6 ^ c8;	// answer: 
		q[2] = c3 ^ c7 ^ c8;
		q[3] = c1 ^ c2 ^ c3 ^ c5 ^ c7 ^ c9;
	end
	
	// the binary expression of the 7-segment display	
	reg[6:0] seg [10:0];
	initial 
	begin
		seg[0] = 7'b0000001;   //  0
		seg[1] = 7'b1001111;   //  1
		seg[2] = 7'b0010010;   //  2
		seg[3] = 7'b0000110;   //  3
		seg[4] = 7'b1001100;   //  4
		seg[5] = 7'b0100100;   //  5
		seg[6] = 7'b0100000;   //  6
		seg[7] = 7'b0001111;   //  7
		seg[8] = 7'b0000000;   //  8
		seg[9] = 7'b0000100;   //  9
		seg[10]= 7'b0111000;   //  F
	end
	
	output wire [6:0] segment_led_1,segment_led_2;
	
	segment timer
	(
		.seg_data_1        (cnt[7:4]),  //seg_data input 
		.seg_data_2        (cnt[3:0]),  //seg_data input 
		.segment_led_1    (segment_led_1),  //MSB~LSB = SEG,DP,G,F,E,D,C,B,A
		.segment_led_2    (segment_led_2)   //MSB~LSB = SEG,DP,G,F,E,D,C,B,A
	);

	always @ (posedge clk) 
	begin
		rd = rd+1; // random value ++ (used for random question)
		fr = fr+1; // count ++ (to stablize the result)
		cd_fr = cd_fr+1; // used for timer count down frequency
		
		if(~btn_fix)  // if btn2 is pressed
		begin
			start = 1; // start the game
			
			// set the timer display
			cnt[7:4] = 4'd3; 
			cnt[3:0] = 4'd0;
			
			lights = q[q_num]; // set LEDs to pre-defined quiz
			
			q_change = 1; // q_change = true, next time use the next question
		end
		
		if(~btn_rand) // if btn0 is pressed
		begin
			start = 1; // start the game
			
			// set the timer display
			cnt[7:4] = 4'd3;
			cnt[3:0] = 4'd0;
			
			// use the current random value (change on every posedge), and try to do xor using the parameters and depending on the random value
			lights = rd[0]*c0 ^ rd[1]*c1 ^ rd[2]*c2 ^ rd[3]*c3 ^ rd[4]*c4 ^ rd[5]*c5 ^ rd[6]*c6 ^ rd[7]*c7 ^ rd[8]*c8 ^ rd[9]*c9;
		end
	
		// if switch changes, set change[x] to "true"
		// Meanwhile, update last[x] (the last state)
		if(sw[9] != last[9])
		begin
			last[9] = sw[9];
			change[9] = 1;	
		end
		if(sw[8] != last[8])
		begin
			last[8] = sw[8];
			change[8] = 1;	
		end
		if(sw[7] != last[7])
		begin
			last[7] = sw[7];
			change[7] = 1;	
		end
		if(sw[6] != last[6])
		begin
			last[6] = sw[6];
			change[6] = 1;	
		end
		if(sw[5] != last[5])
		begin
			last[5] = sw[5];
			change[5] = 1;	
		end
		if(sw[4] != last[4])
		begin
			last[4] = sw[4];
			change[4] = 1;	
		end
		if(sw[3] != last[3])
		begin
			last[3] = sw[3];
			change[3] = 1;	
		end
		if(sw[2] != last[2])
		begin
			last[2] = sw[2];
			change[2] = 1;	
		end
		if(sw[1] != last[1])
		begin
			last[1] = sw[1];
			change[1] = 1;	
		end
		if(sw[0] != last[0])
		begin
			last[0] = sw[0];
			change[0] = 1;	
		end
		
		// xor the lights only when fr == 24'b111111111111111111111111
		// otherwise, it might be "unstable" (prevent over frequent xor operation)
		if(fr == 24'b111111111111111111111111 && start == 1)
		begin
			// Do XOR using the parameters, and depending on whether the switches had been changed during the interval
			lights = lights ^ change[0]*c0 ^ change[1]*c1 ^ change[2]*c2 ^ change[3]*c3 ^ change[4]*c4 ^ change[5]*c5 ^ change[6]*c6 ^ change[7]*c7 ^ change[8]*c8 ^ change[9]*c9;
			change = 10'b0000000000;
			
			// if the lights are all switched off, you win!
			if(lights == 10'b0000000000)
			begin
				// stop the game
				start = 0;
			end
		end
		
		// timer count down only when cd_fr == 26'b11000000000000000000000000
		// this looks like one second on the timer
		if(cd_fr == 26'b11000000000000000000000000 && start == 1)
		begin
			if(cnt[3:0] == 4'd0) 
			begin
				cnt[3:0] = 4'd9; 
				if(cnt[7:4] == 4'd0 ) 
				begin
					cnt[3:0] = 4'd10;
					cnt[7:4] = 4'd10;
				end
				else
				begin
					cnt[7:4] = cnt[7:4] - 1'b1; 
				end
			end
			else cnt[3:0] = cnt[3:0] - 1'b1;
			
			// if time's up, you lose
			if(cnt[3:0] == 4'd10 && cnt[7:4] == 4'd10)
			begin
				// all the lights are switched on
				lights = 10'b1111111111;
				start = 0;
			end
			
			// if q_change == 1 (next question)
			if(q_change == 1)
			begin
				q_num = q_num+1;
				q_change = 0;
			end
			
			// reset cd_fr			
			cd_fr = 26'b00000000000000000000000000;
		end
	end
endmodule

// the module to connect the 7-seg display
module segment
(
input  wire [3:0] seg_data_1,
input  wire [3:0] seg_data_2, 
output wire [6:0] segment_led_1, 
output wire [6:0] segment_led_2  
);
reg[6:0] seg [10:0]; 
initial 
    begin
        seg[0] = 7'b0000001;   //  0
        seg[1] = 7'b1001111;   //  1
        seg[2] = 7'b0010010;   //  2
        seg[3] = 7'b0000110;   //  3
        seg[4] = 7'b1001100;   //  4
        seg[5] = 7'b0100100;   //  5
        seg[6] = 7'b0100000;   //  6
        seg[7] = 7'b0001111;   //  7
        seg[8] = 7'b0000000;   //  8
        seg[9] = 7'b0000100;   //  9
        seg[10]= 7'b0111000;   //  F
    end
   assign segment_led_1 = seg[seg_data_2];
   assign segment_led_2 = seg[seg_data_1];
endmodule 
